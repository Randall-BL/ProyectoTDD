//=======================================================
// ps2.v (con indicador de dato válido)
//=======================================================
module ps2(
    input  wire       iRST_n,
    input  wire       iCLK_50,
    inout  wire       PS2_CLK,
    inout  wire       PS2_DAT,
    output reg [3:0]  char_code,
    output reg        char_valid
);
    // Scancodes...
    localparam SC_0=8'h45, SC_1=8'h16, SC_2=8'h1E, SC_3=8'h26;
    localparam SC_4=8'h25, SC_5=8'h2E, SC_6=8'h36, SC_7=8'h3D;
    localparam SC_8=8'h3E, SC_9=8'h46;
    localparam SC_PLUS=8'h79, SC_MINUS=8'h7B;
    localparam SC_MUL=8'h7C, SC_DIV=8'h4A;
    localparam SC_ENT=8'h5A, SC_BS=8'h66;

    // clk_ps2
    reg [8:0] clk_div;
    wire clk_ps2 = clk_div[8];
    always @(posedge iCLK_50) clk_div<=clk_div+1;

    // sincronización
    reg ps2_clk_i, ps2_clk_d;
    reg ps2_dat_i, ps2_dat_d;
    always @(posedge clk_ps2) begin
        ps2_clk_d<=PS2_CLK; ps2_clk_i<=ps2_clk_d;
        ps2_dat_d<=PS2_DAT; ps2_dat_i<=ps2_dat_d;
    end

    // shift
    reg [10:0] shift;
    reg [3:0]  bit_cnt;
    always @(negedge ps2_clk_i or negedge iRST_n) begin
        if(!iRST_n) begin shift<=0; bit_cnt<=0; end else begin
            shift<= {ps2_dat_i, shift[10:1]};
            bit_cnt<= (bit_cnt==4'd11)?4'd0:bit_cnt+1;
        end
    end

    // decodificación y flag
    always @(posedge clk_ps2 or negedge iRST_n) begin
        if(!iRST_n) begin char_code<=4'hF; char_valid<=0; end
        else if(bit_cnt==4'd11) begin
            char_valid <= 1;
            case(shift[8:1])
                SC_0: char_code<=4'h0; SC_1: char_code<=4'h1;
                SC_2: char_code<=4'h2; SC_3: char_code<=4'h3;
                SC_4: char_code<=4'h4; SC_5: char_code<=4'h5;
                SC_6: char_code<=4'h6; SC_7: char_code<=4'h7;
                SC_8: char_code<=4'h8; SC_9: char_code<=4'h9;
                SC_PLUS:  char_code<=4'hA;
                SC_MINUS: char_code<=4'hB;
                SC_MUL:   char_code<=4'hC;
                SC_DIV:   char_code<=4'hD;
                SC_ENT:   char_code<=4'hE;
                SC_BS:    char_code<=4'hF;
                default:  char_code<=4'hF;
            endcase
        end else char_valid<=0;
    end
endmodule
